module Light_Controller (
    input clk,
    input rst,
    
    // �Է�
    input sw_headlight,      // ���� ������ (SW4)
    input sw_high_beam,      // ����� ����ġ (SW5)
    input [7:0] cds_val,     // ���� ���� ��
    input is_brake,          // �극��ũ
    input turn_left,         // ���� ������
    input turn_right,        // ���� ������
    
    // �� ���: Full Color LED (4�� x 3�� = 12��)
    // [0]:LED1, [1]:LED2, [2]:LED3, [3]:LED4
    output wire [3:0] fc_red,
    output wire [3:0] fc_green,
    output wire [3:0] fc_blue,
    
    // ���: �Ϲ� LED
    output [7:0] led_port
);

    // 1. �������Ʈ �Ǵ�
    wire is_dark = (cds_val < 100); 
    wire head_on = sw_headlight || is_dark; // ������ ON ����
    
    // 2. ������ ���� (White Color: R+G+B ��� ON)
    // ����� (�Ʒ� 2��: LED3, LED4 -> �ε��� 2, 3)
    // ����� (�� 2��: LED1, LED2 -> �ε��� 0, 1)
    
    wire low_beam_on = head_on; 
    wire high_beam_on = head_on && sw_high_beam; // ������ ���� ���¿��� ����� ����ġ

    // ������ LED ���� (Active Low���� High���� Ȯ�� �ʿ�, ���� High=ON)
    // LED 1 (�����)
    assign fc_red[0]   = high_beam_on;
    assign fc_green[0] = high_beam_on;
    assign fc_blue[0]  = high_beam_on;
    
    // LED 2 (�����)
    assign fc_red[1]   = high_beam_on;
    assign fc_green[1] = high_beam_on;
    assign fc_blue[1]  = high_beam_on;
    
    // LED 3 (�����)
    assign fc_red[2]   = low_beam_on;
    assign fc_green[2] = low_beam_on;
    assign fc_blue[2]  = low_beam_on;
    
    // LED 4 (�����)
    assign fc_red[3]   = low_beam_on;
    assign fc_green[3] = low_beam_on;
    assign fc_blue[3]  = low_beam_on;

    // 3. �Ĺ̵�(�̵�/�극��ũ��) PWM (���� ���� ����)
    reg [4:0] pwm_cnt;
    always @(posedge clk) pwm_cnt <= pwm_cnt + 1;
    wire dim_light = pwm_cnt[4]; 
    wire tail_light_on = is_brake ? 1'b1 : (head_on ? dim_light : 1'b0);

    // 4. �Ϲ� LED ���
    assign led_port[7] = turn_left;
    assign led_port[6] = turn_left;
    assign led_port[5] = tail_light_on;
    assign led_port[4] = tail_light_on;
    assign led_port[3] = tail_light_on;
    assign led_port[2] = tail_light_on;
    assign led_port[1] = turn_right;
    assign led_port[0] = turn_right;

endmodule